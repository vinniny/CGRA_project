// ==============================================================================
// CGRA Top-Level Integration - Centralized CSR + Pipelined DMA Architecture
// ==============================================================================
// Integrates:
// - APB CSR interface (control/status registers)
// - Control Unit (3-state FSM with cycle counter)
// - Pipelined DMA Engine (FIFO + separate Read/Write FSMs)
// - CGRA Fabric (4x4 PE array with routing)
// ==============================================================================

module cgra_top #(
    parameter DATA_WIDTH = 32,
    parameter COORD_WIDTH = 4,
    parameter PAYLOAD_WIDTH = 16,
    parameter ADDR_WIDTH = 32,
    parameter SPM_DEPTH = 256,
    parameter RF_DEPTH = 16,
    parameter CONFIG_WIDTH = 64,
    parameter NUM_PES = 16
)(
    input  logic clk,
    input  logic rst_n,
    
    // =========================================================================
    // APB Slave Interface (from CPU/Testbench)
    // =========================================================================
    input  logic                  psel,
    input  logic                  penable,
    input  logic                  pwrite,
    input  logic [ADDR_WIDTH-1:0] paddr,
    input  logic [31:0]           pwdata,
    output logic [31:0]           prdata,
    output logic                  pready,
    output logic                  pslverr,
    
    // =========================================================================
    // AXI4-Lite Master Interface (DMA to External RAM)
    // =========================================================================
    // Write Address Channel
    output logic [ADDR_WIDTH-1:0] m_axi_awaddr,
    output logic                  m_axi_awvalid,
    input  logic                  m_axi_awready,
    
    // Write Data Channel
    output logic [31:0]           m_axi_wdata,
    output logic [3:0]            m_axi_wstrb,
    output logic                  m_axi_wvalid,
    input  logic                  m_axi_wready,
    
    // Write Response Channel
    input  logic                  m_axi_bvalid,
    output logic                  m_axi_bready,
    
    // Read Address Channel
    output logic [ADDR_WIDTH-1:0] m_axi_araddr,
    output logic                  m_axi_arvalid,
    input  logic                  m_axi_arready,
    
    // Read Data Channel
    input  logic [31:0]           m_axi_rdata,
    input  logic                  m_axi_rvalid,
    output logic                  m_axi_rready,
    
    // =========================================================================
    // Interrupt Output
    // =========================================================================
    output logic                  irq,
    
    // =========================================================================
    // Synthesis Keeper (Prevents optimizer from removing unused logic)
    // =========================================================================
    output logic                  synthesis_keep
);

    // =========================================================================
    // Internal Wires: CSR → DMA
    // =========================================================================
    logic [31:0] dma_src;
    logic [31:0] dma_dst;
    logic [31:0] dma_size;
    logic        dma_start;
    logic        dma_busy;
    logic        dma_done;
    
    // =========================================================================
    // Internal Wires: CSR → Control Unit
    // =========================================================================
    logic        cu_start;
    logic        cu_soft_reset;
    logic        cu_busy;
    logic        cu_done;
    logic [31:0] cu_cycles;
    
    // =========================================================================
    // Internal Wires: Control Unit → Array
    // =========================================================================
    logic        pe_enable;
    logic        pe_reset_n;
    logic        array_done;
    
    // =========================================================================
    // Internal Wires: DMA → Tile Memory (Data Fridge)
    // =========================================================================
    logic [11:0] dma_tile_addr;
    logic [1:0]  dma_tile_bank_sel;
    logic        dma_tile_we;
    logic [31:0] dma_tile_wdata;
    logic [31:0] dma_tile_rdata;
    logic        dma_tile_valid;
    
    // Row data from tile memory → Array
    logic [31:0] row_data [0:3];
    logic        row_valid [0:3];
    
    // =========================================================================
    // Internal Wires: DMA → Config Bus (Recipe Book)
    // =========================================================================
    logic [31:0] dma_cfg_addr;
    logic        dma_cfg_we;
    logic [31:0] dma_cfg_wdata;
    logic [3:0]  dma_cfg_pe_sel;  // Which PE to configure (0-15)
    
    // =========================================================================
    // FIX 2: Double-Pump Config Loader (32-bit DMA → 64-bit Config)
    // =========================================================================
    // Protocol: Write High Word (addr[2]=1) → Write Low Word (addr[2]=0) commits 64-bit
    logic [31:0] config_high_reg;     // Holding register for upper 32 bits
    logic [63:0] config_full_word;    // Combined 64-bit config
    logic        config_commit_en;    // Triggers when low word written
    
    always_ff @(posedge clk) begin
        if (!rst_n) begin
            config_high_reg <= 32'd0;
        end else if (dma_cfg_we && dma_cfg_addr[2]) begin
            // Writing to high word address (offset 4 within config slot)
            config_high_reg <= dma_cfg_wdata;
        end
    end
    
    // Commit trigger: DMA writes to low word address (addr[2]=0)
    assign config_commit_en = dma_cfg_we && !dma_cfg_addr[2];
    
    // Combined 64-bit config: {high_reg, current_low_word}
    assign config_full_word = {config_high_reg, dma_cfg_wdata};
    
    // =========================================================================
    // Internal Wires: Control Unit → Flow Control
    // =========================================================================
    logic [3:0]  context_pc;
    logic        global_stall;
    
    // =========================================================================
    // Internal Wires: Configuration (simplified for now)
    // =========================================================================
    logic [CONFIG_WIDTH-1:0] config_frames [0:15];  // 16 PE configs

    // =========================================================================
    // TEMPORARY: Placeholder assignment for config PE selection
    // =========================================================================
    assign dma_cfg_pe_sel = dma_cfg_addr[11:8];  // PE select from higher bits (avoid overlap with slot)
        
    // =========================================================================
    // 1. APB CSR Module
    // =========================================================================
    cgra_apb_csr #(
        .ADDR_WIDTH(ADDR_WIDTH),
        .DATA_WIDTH(32)
    ) u_csr (
        .clk(clk),
        .rst_n(rst_n),
        
        // APB Interface
        .psel(psel),
        .penable(penable),
        .pwrite(pwrite),
        .paddr(paddr),
        .pwdata(pwdata),
        .prdata(prdata),
        .pready(pready),
        .pslverr(pslverr),
        
        // DMA Config Wires
        .dma_src(dma_src),
        .dma_dst(dma_dst),
        .dma_size(dma_size),
        .dma_start(dma_start),
        .dma_busy_i(dma_busy),
        .dma_done_i(dma_done),
        
        // Control Unit Config Wires
        .cu_start(cu_start),
        .cu_soft_reset(cu_soft_reset),
        .cu_busy_i(cu_busy),
        .cu_done_i(cu_done),
        .cu_cycles_i(cu_cycles),
        
        // IRQ
        .irq(irq)
    );
    
    // =========================================================================
    // 2. Pipelined DMA Engine
    // =========================================================================
    cgra_dma_engine #(
        .DATA_WIDTH(32),
        .ADDR_WIDTH(ADDR_WIDTH),
        .FIFO_DEPTH(8)
    ) u_dma (
        .clk(clk),
        .rst_n(rst_n),
        
        // CSR Config
        .cfg_src(dma_src),
        .cfg_dst(dma_dst),
        .cfg_size(dma_size),
        .cfg_start(dma_start),
        .status_busy(dma_busy),
        .status_done(dma_done),
        .irq_done(),  // Not used here - IRQ from CSR
        
        // AXI4-Lite Master
        .m_axi_awaddr(m_axi_awaddr),
        .m_axi_awvalid(m_axi_awvalid),
        .m_axi_awready(m_axi_awready),
        .m_axi_wdata(m_axi_wdata),
        .m_axi_wstrb(m_axi_wstrb),
        .m_axi_wvalid(m_axi_wvalid),
        .m_axi_wready(m_axi_wready),
        .m_axi_bvalid(m_axi_bvalid),
        .m_axi_bready(m_axi_bready),
        .m_axi_araddr(m_axi_araddr),
        .m_axi_arvalid(m_axi_arvalid),
        .m_axi_arready(m_axi_arready),
        .m_axi_rdata(m_axi_rdata),
        .m_axi_rvalid(m_axi_rvalid),
        .m_axi_rready(m_axi_rready),
        
        // Local Memory Interface (To Tile Memory)
        .tile_addr_o(dma_tile_addr),
        .tile_bank_sel_o(dma_tile_bank_sel),
        .tile_we_o(dma_tile_we),
        .tile_wdata_o(dma_tile_wdata),
        
        // Config Interface (To PE Array)
        .config_addr_o(dma_cfg_addr),
        .config_we_o(dma_cfg_we),
        .config_wdata_o(dma_cfg_wdata)
    );
    
    // =========================================================================
    // 3. Control Unit
    // =========================================================================
    cgra_control_unit #(
        .CONTEXT_DEPTH(16),
        .PC_WIDTH(4)
    ) u_cu (
        .clk(clk),
        .rst_n(rst_n),
        
        // CSR Interface
        .start_i(cu_start),
        .soft_reset_i(cu_soft_reset),
        .busy_o(cu_busy),
        .done_o(cu_done),
        .cycle_count_o(cu_cycles),
        
        // Array Interface
        .pe_enable(pe_enable),
        .pe_reset_n(pe_reset_n),
        .array_done_i(array_done),
        
        // Multi-Context Flow Control
        .context_pc_o(context_pc),
        .global_stall_o(global_stall),
        .dma_busy_i(dma_busy),
        
        // Configuration
        .max_cycles_i(32'd0)  // No timeout limit
    );
    
    // =========================================================================
    // 4. Tile Memory (The "Fridge" - Data Banks for PE Array)
    // =========================================================================
    // 4 banks × 1024 words = 16KB total
    // DMA writes to ext_* port, Array reads from bank*_rdata
    cgra_tile_memory #(
        .DATA_WIDTH(DATA_WIDTH),
        .ADDR_WIDTH(12),
        .BANK_DEPTH(1024),
        .NUM_BANKS(4)
    ) u_tile_mem (
        .clk(clk),
        .rst_n(rst_n),
        
        // FIX 3: Dynamic Memory Addressing (Streaming Mode)
        // Each bank address = context_pc, enabling 16-word streaming per run
        
        // Bank 0 (Row 0) - Read port to array
        .bank0_addr({8'd0, context_pc}), // FIX 3: Address = context_pc (0-15)
        .bank0_read(1'b1),               // Always read enabled
        .bank0_write(1'b0),              // Array doesn't write
        .bank0_wdata(32'd0),
        .bank0_rdata(row_data[0]),
        .bank0_valid(row_valid[0]),
        
        // Bank 1 (Row 1) - Read port to array
        .bank1_addr({8'd0, context_pc}), // FIX 3: Address = context_pc
        .bank1_read(1'b1),
        .bank1_write(1'b0),
        .bank1_wdata(32'd0),
        .bank1_rdata(row_data[1]),
        .bank1_valid(row_valid[1]),
        
        // Bank 2 (Row 2) - Read port to array
        .bank2_addr({8'd0, context_pc}), // FIX 3: Address = context_pc
        .bank2_read(1'b1),
        .bank2_write(1'b0),
        .bank2_wdata(32'd0),
        .bank2_rdata(row_data[2]),
        .bank2_valid(row_valid[2]),
        
        // Bank 3 (Row 3) - Read port to array
        .bank3_addr({8'd0, context_pc}), // FIX 3: Address = context_pc
        .bank3_read(1'b1),
        .bank3_write(1'b0),
        .bank3_wdata(32'd0),
        .bank3_rdata(row_data[3]),
        .bank3_valid(row_valid[3]),
        
        // External/DMA port - Write access
        .ext_addr(dma_tile_addr),
        .ext_bank_sel(dma_tile_bank_sel),
        .ext_read(1'b0),             // DMA write only for now
        .ext_write(dma_tile_we),
        .ext_wdata(dma_tile_wdata),
        .ext_rdata(dma_tile_rdata),
        .ext_valid(dma_tile_valid)
    );
    
    // =========================================================================
    // 5. CGRA Array (4x4 PE Mesh)
    // =========================================================================
    
    // =========================================================================
    // AUTO-STOP FEATURE: Programmable Cycle Counter
    // =========================================================================
    // The CPU can program a cycle limit. When the counter reaches 1, array_done
    // is asserted to signal the Control Unit to stop execution automatically.
    //
    // Usage:
    // 1. Write cycle count to cycle_limit register (via CSR or hardcode)
    // 2. Start execution - counter decrements each cycle
    // 3. When counter == 1, array_done pulses to trigger auto-stop
    //
    // For now, we use a simple approach: tie array_done to context_pc overflow
    // This triggers auto-stop after 16 contexts (one complete sweep)
    // More sophisticated: Use a dedicated CSR register for arbitrary counts
    
    // Simple Auto-Stop: Trigger after 16 context cycles (context_pc wraps)
    // This is suitable for single-pass dataflow computations
    logic [4:0] auto_stop_counter;
    logic       auto_stop_armed;
    
    always_ff @(posedge clk) begin
        if (!rst_n) begin
            auto_stop_counter <= 5'd0;
            auto_stop_armed <= 1'b0;
        end else if (cu_soft_reset) begin
            // When CU starts (soft_reset clears then start), arm the counter
            auto_stop_counter <= 5'd0;
            auto_stop_armed <= 1'b1;
        end else if (pe_enable && auto_stop_armed) begin
            // Count while running
            auto_stop_counter <= auto_stop_counter + 1'b1;
        end
    end
    
    // Trigger array_done after 16 cycles (configurable via parameter)
    // This causes the CU to transition to FINISH state
    assign array_done = auto_stop_armed && (auto_stop_counter == 5'd16);
    
    // =========================================================================
    // Edge Output Wires for Synthesis Keeper
    // =========================================================================
    logic [DATA_WIDTH-1:0] edge_n0, edge_n1, edge_n2, edge_n3;
    logic [DATA_WIDTH-1:0] edge_s0, edge_s1, edge_s2, edge_s3;
    logic [DATA_WIDTH-1:0] edge_e0, edge_e1, edge_e2, edge_e3;
    logic [DATA_WIDTH-1:0] edge_w0, edge_w1, edge_w2, edge_w3;
    
    cgra_array_4x4 #(
        .DATA_WIDTH(DATA_WIDTH),
        .COORD_WIDTH(COORD_WIDTH),
        .PAYLOAD_WIDTH(PAYLOAD_WIDTH),
        .ADDR_WIDTH(4),
        .SPM_DEPTH(SPM_DEPTH),
        .RF_DEPTH(RF_DEPTH),
        .CONTEXT_DEPTH(16),
        .PC_WIDTH(4)
    ) u_array (
        .clk(clk),
        .rst_n(rst_n & pe_reset_n),  // Combined reset
        
        // Configuration (simplified - all PEs same config for now)
        .config_frame_00(64'd0),
        .config_frame_01(64'd0),
        .config_frame_02(64'd0),
        .config_frame_03(64'd0),
        .config_frame_10(64'd0),
        .config_frame_11(64'd0),
        .config_frame_12(64'd0),
        .config_frame_13(64'd0),
        .config_frame_20(64'd0),
        .config_frame_21(64'd0),
        .config_frame_22(64'd0),
        .config_frame_23(64'd0),
        .config_frame_30(64'd0),
        .config_frame_31(64'd0),
        .config_frame_32(64'd0),
        .config_frame_33(64'd0),
        .config_valid(1'b0),       // Use config RAM, not direct frame
        
        // Multi-context interface - FIX 2: Double-pump config path
        .context_pc(context_pc),
        .global_stall(global_stall),
        .cfg_wr_addr(dma_cfg_addr[6:3]),         // Config slot address (skip bit 2 used for hi/lo)
        .cfg_wr_data(config_full_word),          // FIX 2: Full 64-bit config
        .cfg_wr_pe_sel(dma_cfg_pe_sel),          // From address decode
        .cfg_wr_en(config_commit_en),            // FIX 2: Only commit on low word write

        
        // North edge inputs - tie off
        .edge_data_in_n0(32'd0),
        .edge_data_in_n1(32'd0),
        .edge_data_in_n2(32'd0),
        .edge_data_in_n3(32'd0),
        .edge_valid_in_n0(1'b0),
        .edge_valid_in_n1(1'b0),
        .edge_valid_in_n2(1'b0),
        .edge_valid_in_n3(1'b0),
        
        // South edge inputs - tie off
        .edge_data_in_s0(32'd0),
        .edge_data_in_s1(32'd0),
        .edge_data_in_s2(32'd0),
        .edge_data_in_s3(32'd0),
        .edge_valid_in_s0(1'b0),
        .edge_valid_in_s1(1'b0),
        .edge_valid_in_s2(1'b0),
        .edge_valid_in_s3(1'b0),
        
        // East edge inputs - tie off
        .edge_data_in_e0(32'd0),
        .edge_data_in_e1(32'd0),
        .edge_data_in_e2(32'd0),
        .edge_data_in_e3(32'd0),
        .edge_valid_in_e0(1'b0),
        .edge_valid_in_e1(1'b0),
        .edge_valid_in_e2(1'b0),
        .edge_valid_in_e3(1'b0),
        
        // West edge inputs - FROM TILE MEMORY (The Data Pipeline!)
        .edge_data_in_w0(row_data[0]),   // Bank 0 -> Row 0 PEs
        .edge_data_in_w1(row_data[1]),   // Bank 1 -> Row 1 PEs
        .edge_data_in_w2(row_data[2]),   // Bank 2 -> Row 2 PEs
        .edge_data_in_w3(row_data[3]),   // Bank 3 -> Row 3 PEs
        .edge_valid_in_w0(row_valid[0]),
        .edge_valid_in_w1(row_valid[1]),
        .edge_valid_in_w2(row_valid[2]),
        .edge_valid_in_w3(row_valid[3]),
        
        // Edge outputs - connected for synthesis keepalive
        .edge_data_out_n0(edge_n0),
        .edge_data_out_n1(edge_n1),
        .edge_data_out_n2(edge_n2),
        .edge_data_out_n3(edge_n3),
        .edge_valid_out_n0(),
        .edge_valid_out_n1(),
        .edge_valid_out_n2(),
        .edge_valid_out_n3(),
        
        .edge_data_out_s0(edge_s0),
        .edge_data_out_s1(edge_s1),
        .edge_data_out_s2(edge_s2),
        .edge_data_out_s3(edge_s3),
        .edge_valid_out_s0(),
        .edge_valid_out_s1(),
        .edge_valid_out_s2(),
        .edge_valid_out_s3(),
        
        .edge_data_out_e0(edge_e0),
        .edge_data_out_e1(edge_e1),
        .edge_data_out_e2(edge_e2),
        .edge_data_out_e3(edge_e3),
        .edge_valid_out_e0(),
        .edge_valid_out_e1(),
        .edge_valid_out_e2(),
        .edge_valid_out_e3(),
        
        .edge_data_out_w0(edge_w0),
        .edge_data_out_w1(edge_w1),
        .edge_data_out_w2(edge_w2),
        .edge_data_out_w3(edge_w3),
        .edge_valid_out_w0(),
        .edge_valid_out_w1(),
        .edge_valid_out_w2(),
        .edge_valid_out_w3()
    );
    
    // =========================================================================
    // Synthesis Keeper: OR-reduce all edge outputs to single bit
    // =========================================================================
    // This prevents the synthesizer from optimizing away the array due to
    // unconnected outputs. Route this pin to a test pad or leave floating.
    assign synthesis_keep = |edge_n0 | |edge_n1 | |edge_n2 | |edge_n3 |
                            |edge_s0 | |edge_s1 | |edge_s2 | |edge_s3 |
                            |edge_e0 | |edge_e1 | |edge_e2 | |edge_e3 |
                            |edge_w0 | |edge_w1 | |edge_w2 | |edge_w3;

endmodule
